Changes made in repo1


hey i am mital

