Changes made in repo1
